
module fadds (
    input  [31:0] fa,
    input  [31:0] fb,
    output [31:0] fres
);
    
endmodule
