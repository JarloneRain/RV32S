

module CPU (
    input clk,
    input rst,
);





endmodule
